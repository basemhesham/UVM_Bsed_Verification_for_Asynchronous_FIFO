package pack1; 
    import uvm_pkg::*;
    `include "uvm_macros.svh"           
    `include "sequence_item.sv"
    `include "sequence.sv"
    `include "sequencer.sv"
    `include "driver.sv"   
    `include "monitor.sv"
    `include "agent.sv"
    `include "subscriber.sv"
    `include "environment.sv"
    `include "test.sv"
endpackage
